--! @file T0_Shutter_Iface_rtl.vhd
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;

library unisim;
use unisim.VComponents.all;

USE work.ipbus.all;

use work.ipbus_reg_types.all;

--! @brief Simple module to generate T0 and shutter signals under IPBus control
--! Similar interface to TPx3_iface_rtl.vhd
--
--! @details
--! \n \n IPBus address map:
--! \li 00 - Activate shutter. Bit 0. Shutter is active if  bit-0=1 , else always 0
--! \li 01 - T0 write to pulse T0. Four cycles of clk_4x ( one cycle of clock sent to DUTs)
--! \li 10 - Delay from signal from accelerator to shutter signal.
--! \li 11 - Which trigger signal to regard as accelerator input. Not currently used.
--! @author David Cussans

entity T0_Shutter_Iface is
  generic (
    g_NUM_ACCELERATOR_SIGNALS: positive := 6 --! Number of hardware signals.
    );
  port (
    clk_4x_i                    : in  std_logic;    --! system clock
    clk_4x_strobe_i               : in  std_logic;    --! strobes high for one cycle every 4 of clk_4x
    accelerator_signals_i       : in std_logic_vector(g_NUM_ACCELERATOR_SIGNALS-1 downto 0); --! hardware signals from accelerator
    T0_o                        : out std_logic;    --! T0 signal retimed onto system clock
    shutter_o                   : out std_logic;    --! shutter signal retimed onto system clock
    ipbus_clk_i                 : IN     std_logic; --! IPBus system clock
    ipbus_i                     : IN     ipb_wbus;
    ipbus_o                     : OUT    ipb_rbus
          
    );     

end entity T0_Shutter_Iface;

architecture rtl of T0_Shutter_Iface is

  signal s_T0 , s_T0_d1 , s_T0_d2 , s_stretch_T0_in: std_logic := '0';  --! signal after IBufDS and sampled onto clk_4x
  signal s_stretch_T0_in_sr : std_logic_vector(2 downto 0) := "111"; --! Gets shifted out by clk_4x logic. Loaded by T0ger_i
  signal s_T0_out_sr : std_logic_vector(2 downto 0) := "111"; --! Gets shifted out by clk_4x logic. Loaded by strobe_4x_logic

  signal s_shutter , s_shutter_d1 , s_shutter_d2 : std_logic := '0';  --! signal after IBufDS and sampled onto clk_4x
  signal s_shutter_delay : std_logic_vector(ipbus_i.ipb_wdata'range); --! 
  signal s_T0_ipbus , s_T0_ipbus_d1 , s_T0_ipbus_d2: std_logic := '0';  --! T0 sync signal
  signal s_shutter_ipbus , s_shutter_ipbus_d1 , s_shutter_ipbus_d2 , s_shutter_ipbus_enable: std_logic := '0';  -- Signals that get combined with incoming hardware signals from TPIx3 telescope
  signal s_accelerator_trigger_shutter : std_logic := '0'; --! Taking this line high triggers a shutter
                                                                             
  signal s_ipbus_ack      : std_logic := '0';  -- used to produce a delayed IPBus ack signal
  signal s_counting_down  : std_logic ; -- high whilst counting down then goes low.
  
begin  -- architecture rtl

  --------------------
    ipbus_write: process (ipbus_clk_i)
    begin  -- process ipb_clk_i
    if rising_edge(ipbus_clk_i) then
        s_T0_ipbus <= '0';
        if (ipbus_i.ipb_strobe = '1' and ipbus_i.ipb_write = '1') then
            case ipbus_i.ipb_addr(1 downto 0) is
              when "00" => s_shutter_ipbus_enable <= ipbus_i.ipb_wdata(0) ; -- Set IPBus shutter enable
              when "01" => s_T0_ipbus <= '1'; -- set T0 signal high
              when "10" => s_shutter_delay <= ipbus_i.ipb_wdata;
              when others => null;
            end case;
        end if;
        s_ipbus_ack <= ipbus_i.ipb_strobe and not s_ipbus_ack;
    end if;
    end process ipbus_write;

    ipbus_o.ipb_ack <= s_ipbus_ack;
    ipbus_o.ipb_err <= '0';


    ------------------
    -- Bodge - just wire up trigger input 5 to the accelerator signal for now.
    s_accelerator_trigger_shutter <= accelerator_signals_i(g_NUM_ACCELERATOR_SIGNALS-1);

    cmp_delayPulse: entity work.DelayPulse4x
      generic map (
        g_MAX_WIDTH => s_shutter_delay'length )
    port map (
      clk_4x_i          => clk_4x_i,
      clk_4x_strobe_i   => clk_4x_strobe_i,
      delay_cycles_i    => s_shutter_delay,
      pulse_i           => s_accelerator_trigger_shutter,
      pulse_o           => shutter_o
      );


    --! Retime T0 generated by IPBus onto clk_4x and align with strobe
    cmp_T0_retime: entity work.stretchPulse4x
      port map (
        clk_4x_i      => clk_4x_i,
        clk_4x_strobe_i => clk_4x_strobe_i,
        pulse_i       => s_T0_ipbus,
        pulse_o       => T0_o);

    

end architecture rtl;
